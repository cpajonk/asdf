module asdf

const myconst = 'myconst'

pub fn do_thing() {
	println(asdf.myconst)
}

fn do_internal_thing() int {
	return 10
}
