module asdf

const myconst = 'myconst'

pub fn do_thing() {
	println(asdf.myconst)
}
